** Fractional Order Sallen Key LPF - Winter Training (30/EC/14)

.lib eval.lib

** Fractional Capacitance Simulation - Order = 1.5 C(Beta)
Rax 3 200 111.1
Rbx 200 300 251.7
Rcx 300 400 378.7
Rdx 400 500 888.9
Rex 500 0 7.369k
Cbx 200 300 83.8nF
Ccx 300 400 0.296uF
Cdx 400 500 0.537uF
Cex 500 0 0.695uF

** Fractional Capacitance Simulation - Order = 1.1 C(Alpha)
Ray 2 20 658.7
Rby 20 30 196.3
Rcy 30 40 134.6
Rdy 40 50 159.0
Rey 50 6 369.5
Cby 20 30 68.9nF
Ccy 30 40 0.627uF
Cdy 40 50 2.18uF
Cey 50 6 6.64uF

** Sallen Key Ckt
R1 1 2 1k
R2 2 3 2k
R3 4 0 3k
R4 4 6 4k
X1 3 4 71 41 6 UA741
Vcc+ 71 0 dc 12V
Vcc- 41 0 dc -12V
Vin 1 0 ac 1V

.ac dec 50 1Hz 1MegHz
.probe
.end