** Fractional Order KHN simulation - Winter Training (30/EC/14)

.lib eval.lib

** Fractional Capacitance Simulation - Order = 1.5 C(alpha)
Rax 7 200 111.1
Rbx 200 300 251.7
Rcx 300 400 378.7
Rdx 400 500 888.9
Rex 500 8 7.369k
Cbx 200 300 83.8nF
Ccx 300 400 0.296uF
Cdx 400 500 0.537uF
Cex 500 8 0.695uF

** Fractional Capacitance Simulation - Order = 1.1 C(Beta)
Ray 5 20 658.7
Rby 20 30 196.3
Rcy 30 40 134.6
Rdy 40 50 159.0
Rey 50 6 369.5
Cby 20 30 68.9nF
Ccy 30 40 0.627uF
Cdy 40 50 2.18uF
Cey 50 6 6.64uF

** KHN Ckt
X1 2 3 71 41 4 UA741
X2 0 5 72 42 6 UA741
X3 0 7 73 43 8 UA741
R1 4 5 1k
R2 6 7 2k
R3 2 6 3k
R4 1 2 4k
R5 3 4 5k
R6 3 8 6k
Vcc1+ 71 0 dc 12V
Vcc1- 41 0 dc -12V
Vcc2+ 72 0 dc 12V
Vcc2- 42 0 dc -12V
Vcc3+ 73 0 dc 12V
Vcc3- 43 0 dc -12V
Vin 1 0 ac 1V

.ac dec 50 1Hz 1MegHz
.probe
.end